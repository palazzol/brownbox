.title KiCad schematic

X1 Vcc GNDREF PowerIn

R1 A VCC 2K
R4 Net-_D1-Pad2_ GNDREF 2K
R6 Net-_C2-Pad1_ GNDREF 220K
C1 Net-_C1-Pad1_ Net-_C1-Pad2_ 390pF
C2 Net-_C2-Pad1_ Net-_C2-Pad2_ 330pF
R3 Net-_D1-Pad2_ Net-_C1-Pad2_ 2K
R2 Net-_C2-Pad2_ A 2K
Q1 GNDREF Net-_C1-Pad1_ A 2N5134
RV1 VCC Net-_R5-Pad1_ Net-_R5-Pad1_ 100K
Q2 VCC Net-_C2-Pad1_ Net-_D1-Pad2_ 2N5139
R5 Net-_R5-Pad1_ Net-_C1-Pad1_ 150K

R7 B VCC 2K
R10 S11C2 GNDREF 2K
R12 Net-_C4-Pad1_ GNDREF 220K
C3 Net-_C3-Pad1_ Net-_C3-Pad2_ 0.1uF
C4 Net-_C4-Pad1_ Net-_C4-Pad2_ 0.2uF
R9 S11C2 Net-_C3-Pad2_ 2K
R8 Net-_C4-Pad2_ B 2K
Q3 GNDREF Net-_C3-Pad1_ B 2N5134
RV2 VCC Net-_R11-Pad1_ Net-_R11-Pad1_ 100K
R11 Net-_R11-Pad1_ Net-_C3-Pad1_ 150K
Q4 VCC Net-_C4-Pad1_ S11C2 2N5139

.end